`timescale 1ns/1ns
module part1_tb();

logic [31:0] X, Y, out;

part1 DUT(X, Y, out);

initial begin

	X = 32'b00000000000000000000000000000000;
	Y = 32'b00000000000000000000000000000000;
	
	#10;
	
	X = 32'b1100_0001_1001_0000_0000_0000_0000_0000;
	Y = 32'b0100_0001_0001_1000_0000_0000_0000_0000;
	
	#10;
	
	$stop();
	
end

endmodule
