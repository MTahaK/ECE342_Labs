`timescale 1ns/1ns
module part2tb();

logic [16:0] X, Y, result;
logic [22:0] X_22, Y_22, result_22;
logic [24:0] X_24, Y_24, result_24;
// logic [64:0] X_64, Y_64, result_64;
wire zero, underflow, overflow, nan;
wire zero_22, underflow_22, overflow_22, nan_22;
wire zero_24, underflow_24, overflow_24, nan_24;


part2 DUT(X, Y, result, zero, underflow, overflow, nan);
defparam DUT.M = 8;
defparam DUT.E = 8;
part2 DUT_22(X_22, Y_22, result_22, zero_22, underflow_22, overflow_22,nan_22);
defparam DUT_22.M = 16;
defparam DUT_22.E = 6;
part2 DUT_24(X_24, Y_24, result_24, zero_24, underflow_24, overflow_24, nan_24);
defparam DUT_24.M = 8;
defparam DUT_24.E = 16;
// part2 DUT64(X_64, Y_64, result_64, zero_64, underflow_64, overflow_64, nan_64);
// defparam DUT64.E = 11;
// defparam DUT64.M = 52;


initial begin

	
	
	

    // #5;

    // X = 'h1d0bc;
    // Y = 'h1a67a;
	// // X_64 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    // // Y_64 = 64'b0000000000000000000000000000000000000000000000000000000000000000;


    // #5;

    

    // #5;

    // // X = 32'b1100_0001_1001_0000_0000_0000_0000_0000;
    // // Y = 32'b0100_0001_0001_1000_0000_0000_0000_0000;
	// X_22 = 'h1f08a3;
	// Y_22 = 'h3f0001;
	// // X_64 = 64'b1100_0001_1001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    // // Y_64 = 64'b0100_0001_0001_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
	

    // // Result = 1100_0011_0010_1011_0000_0000_0000_0000

    // #5;


    // #5;

    //Zero case
    // X = 32'b1000_0000_0000_0000_0000_0000_0000_0000; // E = 0, M = 0
    // Y = 32'b0100_0001_0001_1111_0110_0000_0000_0000;
	X_24 = 'h11bf838;
	Y_24 = 'h199e402;
	// X_64 = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    // Y_64 = 64'b0100_0001_0001_1111_0110_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

    #5;

    

    #5;

    //Underflow case
    // X = 32'b1000_1111_0000_0000_1111_1111_0000_0000; //E = 30
    // Y = 32'b0001_0100_0001_1000_0000_0000_1111_1111; //E = 40
	X_24 = 'h0fffd01;
	Y_24 = 'h0fffd01;
	// X_64 = 64'b1000_1111_0000_0000_1111_1111_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    // Y_64 = 64'b0001_0100_0001_1000_0000_0000_1111_1111_0000_0000_0000_0000_0000_0000_0000_0000;

    #5;

    // #5;

    // //Not-a-Number case
    // // X = 32'b1000_0000_0000_0000_0000_0000_0000_0000; // Zero
    // // Y = 32'b0111_1111_1000_0000_0000_0000_0000_0000; // Infinity
	// // X_64 = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    // // Y_64 = 64'b0111_1111_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

    // #5;

   

    // #5;

    // //Overflow case
    // // X = 32'b1111_1111_1000_0000_1111_1111_0000_0000; //E = 256
    // // Y = 32'b0111_1111_1001_1000_0000_0000_1111_1111; //E = 256
	// X_64 = 64'b1111_1111_1000_0000_1111_1111_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    // Y_64 = 64'b0111_1111_1001_1000_0000_0000_1111_1111_0000_0000_0000_0000_0000_0000_0000_0000;

    #5;
    $stop();
	
end

endmodule
