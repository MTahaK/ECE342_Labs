module wallace_mult #(width=8) (
    input [7:0] x,
    input [7:0] y,
    output [15:0] out  	
);

// Wires corresponding to each level of the WTM. 
wire [15:0] s_lev[0:3][1:2];
wire [15:0] c_lev[0:3][1:2];

// Rest of your code goes here. 


endmodule


