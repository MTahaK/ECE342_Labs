
module nios_system (
	clk_clk);	

	input		clk_clk;
endmodule
